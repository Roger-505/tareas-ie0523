module tester_parkingController(
     output         vehicle_arrival
    ,output [ 15:0] code
    ,output         vehicle_left  
    ,output    clk
    ,output    rst
);

endmodule

`ifndef STATE_DEFS_VH
`define STATE_DEFS_VH

`define NO_VEHICLE      6'd  1
`define WAIT_FOR_PIN    6'd  2
`define INCORRECT_PIN   6'd  4
`define CORRECT_PIN     6'd  8
`define WAIT_TO_CLOSE   6'd 16
`define BLOCKED         6'd 32
`define DEFAULT         6'd  0

`endif
